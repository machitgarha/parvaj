library ieee;
use ieee.std_logic_1164.all;

entity <entity-name> is
end entity;

architecture <architecture-name> of <entity-name> is
<component>
begin
    instance: <source-entity-name> port map(

    );
end architecture;
