library ieee;
use ieee.std_logic_1164.all;

entity <entity-name> is
    port(

    );
end entity;

architecture <architecture-name> of <entity-name> is
begin

end architecture;
